module full_adder(sum, cout, a, b, cin);
    output sum, cout;
    input  a, b, cin;
    wire   partial_s, partial_c1, partial_c2;

    xor x0(partial_s, a, b);
    xor x1(sum, partial_s, cin);
    and a0(partial_c1, a, b);
    and a1(partial_c2, partial_s, cin);
    or  o1(cout, partial_c1, partial_c2);
endmodule // full_adder


`define ALU_ADD    3'h2
`define ALU_SUB    3'h3
`define ALU_AND    3'h4
`define ALU_OR     3'h5
`define ALU_NOR    3'h6
`define ALU_XOR    3'h7

// 01x -> arithmetic, 1xx -> logic
module alu1(out, carryout, A, B, carryin, control);
    output      out, carryout;
    input       A, B, carryin;
    input [2:0] control;
    // add code here!!!
	wire wad, wsb, warith, wlog, couta, couts, cout1, cout2, Bin;
	
	not n0(Bin, B);
	full_adder ad1(wad, couta, A, B, carryin);
	full_adder sb1(wsb, couts, A, Bin, carryin);
	mux2 m0(warith, wad, wsb, control[0]);
	mux2 m1(cout1, couta, couts, control[0]);
	logicunit l0(wlog, A, B, control[1:0]);
	mux2 m2(out, warith, wlog, control[2]);	
	assign cout2 = 1'h0;
	mux2 m3(carryout, cout1, cout2, control[2]);
	

endmodule // alu1
